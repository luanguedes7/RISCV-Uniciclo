
library ieee ;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

entity control is
    port (
	opcode : in std_logic_vector(6 downto 0);
	func3 : in std_logic_vector(2 downto 0);
	branch : out std_logic;
	mem_read : out std_logic;
	mem_to_reg : out std_logic;
	alu_op : out std_logic_vector(1 downto 0);
	mem_write : out std_logic;
	alu_src: out std_logic;
	reg_write: out std_logic;
	reg_write_src : out std_logic_vector(1 downto 0);
	mem_byte_en : out std_logic;
	mem_sgn_en : out std_logic
    );
end control;

architecture arc of control is
begin
    process (opcode) is
    begin
	case opcode is
	    when "0110011" => -- R type
		branch <= '0';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "11";
		mem_write <= '0';
		alu_src <= '0';
		reg_write <= '1';
		reg_write_src <= "00";
		mem_byte_en <= '0';
		mem_sgn_en <= '0';
	    when "0010011" => -- I type (logic)
		branch <= '0';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "10";
		mem_write <= '0';
		alu_src <= '1';
		reg_write <= '1';
		reg_write_src <= "00";
		mem_byte_en <= '0';
		mem_sgn_en <= '0';
	    when "0000011" => -- I type (load)
		branch <= '0';
		mem_read <= '1';
		mem_to_reg <= '1';
		alu_op <= "00";
		mem_write <= '0';
		alu_src <= '1';
		reg_write <= '1';
		reg_write_src <= "00";
		
		if func3(1 downto 0) = "00" then
		    mem_byte_en <= '1';
		else
		    mem_byte_en <= '0';
		end if;
		if func3 = "100" then
		    mem_sgn_en <= '1';
		else
		    mem_sgn_en <= '0';
		end if;
	    when "1100111" => -- I type (jaur)
		branch <= '1';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "00";
		mem_write <= '0';
		alu_src <= '1';
		reg_write <= '1';
		reg_write_src <= "11";
		mem_byte_en <= '0';
		mem_sgn_en <= '0';
	    when "0100011" => -- S type
		branch <= '0';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "00";
		mem_write <= '1';
		alu_src <= '1';
		reg_write <= '0';
		reg_write_src <= "00";
		if func3 = "000" then
		    mem_byte_en <= '1';
		else
		    mem_byte_en <= '0';
		end if;
		mem_sgn_en <= '0';
	    when "1100011" => -- SB type
		branch <= '1';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "01";
		mem_write <= '0';
		alu_src <= '0';
		reg_write <= '0';
		reg_write_src <= "00";
		mem_byte_en <= '0';
		mem_sgn_en <= '0';
	    when "0110111" => -- U type (lui)
		branch <= '0';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "00";
		mem_write <= '0';
		alu_src <= '0';
		reg_write <= '1';
		reg_write_src <= "01";
		mem_byte_en <= '0';
		mem_sgn_en <= '0';
	    when "0010111" => -- U type (aiupc)
		branch <= '0';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "00";
		mem_write <= '0';
		alu_src <= '0';
		reg_write <= '1';
		reg_write_src <= "10";
		mem_byte_en <= '0';
		mem_sgn_en <= '0';
	    when "1101111" => -- UJ type (jal)
		branch <= '1';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "00";
		mem_write <= '0';
		alu_src <= '1';
		reg_write <= '1';
		reg_write_src <= "11";
		mem_byte_en <= '0';
		mem_sgn_en <= '0';
	when others =>
		branch <= '0';
		mem_read <= '0';
		mem_to_reg <= '0';
		alu_op <= "00";
		mem_write <= '0';
		alu_src <= '0';
		reg_write <= '0';
		reg_write_src <= "00";
		mem_byte_en <= '0';
		mem_sgn_en <= '0';
	end case;
    end process;

end arc;



library ieee ;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use std.textio.all;

entity unicycle_riscv_tb is
end unicycle_riscv_tb;

architecture tb of unicycle_riscv_tb is
    signal clk : std_logic := '0';
    constant clk_period : time := 10 ns;
    signal rst : std_logic := '1';
    component unicycle_riscv is
	port (
	    clk : in std_logic;
	    pc_rst : in std_logic
   	);
    end component;

begin
    process is
    begin
        clk <= '1';
        wait for clk_period / 2;
        clk <= '0';
        wait for clk_period / 2;
	if (rst = '1') then rst <= '0'; end if;
    end process;
    
    dut : unicycle_riscv
    port map (
	clk => clk,
	pc_rst => rst
    );

    process is
	variable i : integer;
	file text_file: TEXT open read_mode is "code.asm";
	variable text_line: line;
	variable str : string(1 to 100);
	variable size : natural;
    begin
	readline(text_file, text_line);
	while not endfile(text_file) loop
	    readline(text_file, text_line);
	    if text_line'length > 0 then
		str := (others => ' ');
		read(text_line, str(1 to text_line'length));

		report str;
	    end if;
	    wait for clk_period;
	end loop;
	wait;
    end process;

end tb;